* C:\Users\felipe\Desktop\DEV\Circuitos El�tricos\Lab3\Lab3-6-v2.sch

* Schematics Version 9.1 - Web Update 1
* Wed May 22 19:29:52 2024



** Analysis setup **
.tran 0ns 1ms 0 1us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Lab3-6-v2.net"
.INC "Lab3-6-v2.als"


.probe


.END
