* C:\Users\felipe\Desktop\DEV\Circuitos El�tricos\Lab2\Lab2-4.sch

* Schematics Version 9.1 - Web Update 1
* Tue Apr 23 18:44:33 2024



** Analysis setup **
.ac DEC 10 10Hz 1GHz
.tran 0us 20ms 0 10u
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Lab2-4.net"
.INC "Lab2-4.als"


.probe


.END
