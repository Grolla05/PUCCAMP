* C:\Users\felipe\Desktop\DEV\Circuitos El�tricos\Lab4\Amostrador-FPB-Final.sch

* Schematics Version 9.1 - Web Update 1
* Wed May 29 08:25:56 2024



** Analysis setup **
.tran 0s 10ms 0 10us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Amostrador-FPB-Final.net"
.INC "Amostrador-FPB-Final.als"


.probe


.END
