* C:\Users\felipe\Desktop\DEV\Circuitos El�tricos\Lab4\Cod-Prioridade-Final.sch

* Schematics Version 9.1 - Web Update 1
* Wed May 29 18:01:24 2024



** Analysis setup **
.tran 0 10ms 0 1ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Cod-Prioridade-Final.net"
.INC "Cod-Prioridade-Final.als"


.probe


.END
