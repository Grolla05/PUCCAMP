* C:\Users\felipe\Desktop\DEV\Circuitos El�tricos\Lab3\Lab3-8-v2.sch

* Schematics Version 9.1 - Web Update 1
* Tue May 21 18:44:04 2024



** Analysis setup **
.tran 0ns 1ms 0 1us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Lab3-8-v2.net"
.INC "Lab3-8-v2.als"


.probe


.END
