* C:\Users\felipe\Desktop\Eletronica\Senoide_Cap.sch

* Schematics Version 9.1 - Web Update 1
* Tue Mar 19 20:42:47 2024



** Analysis setup **
.tran 0s 16.67ms 0 10us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Senoide_Cap.net"
.INC "Senoide_Cap.als"


.probe


.END
