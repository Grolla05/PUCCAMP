* C:\Users\felipe\Desktop\DEV\Circuitos El�tricos\Circuito 1.sch

* Schematics Version 9.1 - Web Update 1
* Mon Feb 26 20:48:22 2024



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Circuito 1.net"
.INC "Circuito 1.als"


.probe


.END
