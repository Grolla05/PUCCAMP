* C:\Users\felipe\Desktop\DEV\Circuitos El�tricos\LAB1\Lab 1-1-1.sch

* Schematics Version 9.1 - Web Update 1
* Thu Mar 28 16:25:27 2024



** Analysis setup **
.tran 0s 100ms 0 10us
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Lab 1-1-1.net"
.INC "Lab 1-1-1.als"


.probe


.END
